module fir_57tap_lowpass (
    input  wire              clk,
    input  wire signed [15:0] data_in,
    output reg  signed [15:0] data_out
);

    // Hệ số FIR (fixed point Q1.14, nhân với 16384)
    reg signed [15:0] coeffs [0:56];
    initial begin
   coeffs[0]   = -3;    // -0.000164 * 16384
       coeffs[0] = -1; // -0.000085 * 16384
coeffs[1] = -2; // -0.000098 * 16384
coeffs[2] = -1; // -0.000076 * 16384
coeffs[3] = 0; // 0.000000 * 16384
coeffs[4] = 3; // 0.000154 * 16384
coeffs[5] = 7; // 0.000411 * 16384
coeffs[6] = 13; // 0.000799 * 16384
coeffs[7] = 22; // 0.001345 * 16384
coeffs[8] = 34; // 0.002076 * 16384
coeffs[9] = 49; // 0.003016 * 16384
coeffs[10] = 69; // 0.004184 * 16384
coeffs[11] = 92; // 0.005595 * 16384
coeffs[12] = 119; // 0.007255 * 16384
coeffs[13] = 150; // 0.009162 * 16384
coeffs[14] = 185; // 0.011303 * 16384
coeffs[15] = 224; // 0.013657 * 16384
coeffs[16] = 265; // 0.016190 * 16384
coeffs[17] = 309; // 0.018862 * 16384
coeffs[18] = 354; // 0.021618 * 16384
coeffs[19] = 400; // 0.024401 * 16384
coeffs[20] = 445; // 0.027146 * 16384
coeffs[21] = 488; // 0.029784 * 16384
coeffs[22] = 528; // 0.032245 * 16384
coeffs[23] = 565; // 0.034463 * 16384
coeffs[24] = 596; // 0.036375 * 16384
coeffs[25] = 621; // 0.037924 * 16384
coeffs[26] = 640; // 0.039066 * 16384
coeffs[27] = 652; // 0.039765 * 16384
coeffs[28] = 655; // 0.040000 * 16384
coeffs[29] = 652; // 0.039765 * 16384
coeffs[30] = 640; // 0.039066 * 16384
coeffs[31] = 621; // 0.037924 * 16384
coeffs[32] = 596; // 0.036375 * 16384
coeffs[33] = 565; // 0.034463 * 16384
coeffs[34] = 528; // 0.032245 * 16384
coeffs[35] = 488; // 0.029784 * 16384
coeffs[36] = 445; // 0.027146 * 16384
coeffs[37] = 400; // 0.024401 * 16384
coeffs[38] = 354; // 0.021618 * 16384
coeffs[39] = 309; // 0.018862 * 16384
coeffs[40] = 265; // 0.016190 * 16384
coeffs[41] = 224; // 0.013657 * 16384
coeffs[42] = 185; // 0.011303 * 16384
coeffs[43] = 150; // 0.009162 * 16384
coeffs[44] = 119; // 0.007255 * 16384
coeffs[45] = 92; // 0.005595 * 16384
coeffs[46] = 69; // 0.004184 * 16384
coeffs[47] = 49; // 0.003016 * 16384
coeffs[48] = 34; // 0.002076 * 16384
coeffs[49] = 22; // 0.001345 * 16384
coeffs[50] = 13; // 0.000799 * 16384
coeffs[51] = 7; // 0.000411 * 16384
coeffs[52] = 3; // 0.000154 * 16384
coeffs[53] = 0; // 0.000000 * 16384
coeffs[54] = -1; // -0.000076 * 16384
coeffs[55] = -2; // -0.000098 * 16384
coeffs[56] = -1; // -0.000085 * 16384

    end

    // Dãy giá trị đầu vào
    reg signed [15:0] x_reg [0:56];

    // Cập nhật dãy mẫu vào và tính toán kết quả
    integer i;
    reg signed [31:0] acc;

    always @(posedge clk) begin
        // Dịch mẫu vào
        for (i = 56; i > 0; i = i - 1)
            x_reg[i] <= x_reg[i - 1];
        x_reg[0] <= data_in;

        // Tính tích chập (convolution)
        acc = 0;
        for (i = 0; i < 57; i = i + 1)
            acc = acc + x_reg[i] * coeffs[i];

        // Chia lại độ lớn nếu cần (ví dụ >>14 cho hệ số Q1.14)
        data_out <= acc >>> 14;
    end

endmodule
