module fir_57tap_bandpass (
    input  wire              clk,
    input  wire signed [15:0] data_in,
    output reg  signed [15:0] data_out
);

    // Hệ số FIR (fixed-point Q1.14, nhân với 16384)
    reg signed [15:0] coeffs [0:56];
    initial begin
           coeffs[0]  = -1;    // -0.000078 * 16384
    coeffs[1]  = -2;    // -0.000144 * 16384
    coeffs[2]  = -3;    // -0.000153 * 16384
    coeffs[3]  = 0;     // -0.000000 * 16384
    coeffs[4]  = 7;     // 0.000447 * 16384
    coeffs[5]  = 21;    // 0.001301 * 16384
    coeffs[6]  = 43;    // 0.002611 * 16384
    coeffs[7]  = 70;    // 0.004297 * 16384
    coeffs[8]  = 100;   // 0.006118 * 16384
    coeffs[9]  = 125;   // 0.007656 * 16384
    coeffs[10] = 137;   // 0.008357 * 16384
    coeffs[11] = 125;   // 0.007620 * 16384
    coeffs[12] = 81;    // 0.004928 * 16384
    coeffs[13] = 0;     // 0.000000 * 16384
    coeffs[14] = -116;  // -0.007073 * 16384
    coeffs[15] = -257;  // -0.015735 * 16384
    coeffs[16] = -409;  // -0.024964 * 16384
    coeffs[17] = -546;  // -0.033366 * 16384
    coeffs[18] = -644;  // -0.039371 * 16384
    coeffs[19] = -678;  // -0.041499 * 16384
    coeffs[20] = -633;  // -0.038659 * 16384
    coeffs[21] = -498;  // -0.030406 * 16384
    coeffs[22] = -280;  // -0.017112 * 16384
    coeffs[23] = 0;     // 0.000000 * 16384
    coeffs[24] = 311;   // 0.018980 * 16384
    coeffs[25] = 613;   // 0.037424 * 16384
    coeffs[26] = 865;   // 0.052845 * 16384
    coeffs[27] = 1032;  // 0.063081 * 16384
    coeffs[28] = 1093;  // 0.066667 * 16384
    coeffs[29] = 1032;  // 0.063081 * 16384
    coeffs[30] = 865;   // 0.052845 * 16384
    coeffs[31] = 613;   // 0.037424 * 16384
    coeffs[32] = 311;   // 0.018980 * 16384
    coeffs[33] = 0;     // 0.000000 * 16384
    coeffs[34] = -280;  // -0.017112 * 16384
    coeffs[35] = -498;  // -0.030406 * 16384
    coeffs[36] = -633;  // -0.038659 * 16384
    coeffs[37] = -678;  // -0.041499 * 16384
    coeffs[38] = -644;  // -0.039371 * 16384
    coeffs[39] = -546;  // -0.033366 * 16384
    coeffs[40] = -409;  // -0.024964 * 16384
    coeffs[41] = -257;  // -0.015735 * 16384
    coeffs[42] = -116;  // -0.007073 * 16384
    coeffs[43] = 0;     // -0.000000 * 16384
    coeffs[44] = 81;    // 0.004928 * 16384
    coeffs[45] = 125;   // 0.007620 * 16384
    coeffs[46] = 137;   // 0.008357 * 16384
    coeffs[47] = 125;   // 0.007656 * 16384
    coeffs[48] = 100;   // 0.006118 * 16384
    coeffs[49] = 70;    // 0.004297 * 16384
    coeffs[50] = 43;    // 0.002611 * 16384
    coeffs[51] = 21;    // 0.001301 * 16384
    coeffs[52] = 7;     // 0.000447 * 16384
    coeffs[53] = 0;     // -0.000000 * 16384
    coeffs[54] = -3;    // -0.000153 * 16384
    coeffs[55] = -2;    // -0.000144 * 16384
    coeffs[56] = -1;    // -0.000078 * 16384

    end

    // Dãy mẫu đầu vào
    reg signed [15:0] x_reg [0:56];

    // Biến dùng trong xử lý
    integer i;
    reg signed [31:0] acc;

    always @(posedge clk) begin
        // Dịch dữ liệu
        for (i = 56; i > 0; i = i - 1)
            x_reg[i] <= x_reg[i - 1];
        x_reg[0] <= data_in;

        // Tính tích chập
        acc = 0;
        for (i = 0; i < 57; i = i + 1)
            acc = acc + x_reg[i] * coeffs[i];

        // Chia lại độ lớn (chuẩn Q1.14)
        data_out <= acc >>> 14;
    end

endmodule
