module fir_57tap_highpass (
    input  wire              clk,
    input  wire signed [15:0] data_in,
    output reg  signed [15:0] data_out
);

    // Hệ số FIR (fixed-point Q1.14, nhân với 16384)
    reg signed [15:0] coeffs [0:56];
    initial begin
            coeffs[0]  = 0;     // 0.000024 * 16384
    coeffs[1]  = 3;     // 0.000206 * 16384
    coeffs[2]  = 8;     // 0.000511 * 16384
    coeffs[3]  = 14;    // 0.000877 * 16384
    coeffs[4]  = 19;    // 0.001169 * 16384
    coeffs[5]  = 20;    // 0.001200 * 16384
    coeffs[6]  = 13;    // 0.000778 * 16384
    coeffs[7]  = -4;    // -0.000219 * 16384
    coeffs[8]  = -29;   // -0.001766 * 16384
    coeffs[9]  = -60;   // -0.003631 * 16384
    coeffs[10] = -88;   // -0.005364 * 16384
    coeffs[11] = -104;  // -0.006354 * 16384
    coeffs[12] = -98;   // -0.005959 * 16384
    coeffs[13] = -60;   // -0.003686 * 16384
    coeffs[14] = 10;    // 0.000602 * 16384
    coeffs[15] = 107;   // 0.006529 * 16384
    coeffs[16] = 215;   // 0.013124 * 16384
    coeffs[17] = 309;   // 0.018880 * 16384
    coeffs[18] = 360;   // 0.021956 * 16384
    coeffs[19] = 336;   // 0.020507 * 16384
    coeffs[20] = 214;   // 0.013077 * 16384
    coeffs[21] = -17;   // -0.001012 * 16384
    coeffs[22] = -350;  // -0.021385 * 16384
    coeffs[23] = -761;  // -0.046516 * 16384
    coeffs[24] = -1209; // -0.073855 * 16384
    coeffs[25] = -1641; // -0.100173 * 16384
    coeffs[26] = -1999; // -0.122078 * 16384
    coeffs[27] = -2238; // -0.136589 * 16384
    coeffs[28] = 14060661; // 0.858333 * 16384
    coeffs[29] = -2238; // -0.136589 * 16384
    coeffs[30] = -1999; // -0.122078 * 16384
    coeffs[31] = -1641; // -0.100173 * 16384
    coeffs[32] = -1209; // -0.073855 * 16384
    coeffs[33] = -761;  // -0.046516 * 16384
    coeffs[34] = -350;  // -0.021385 * 16384
    coeffs[35] = -17;   // -0.001012 * 16384
    coeffs[36] = 214;   // 0.013077 * 16384
    coeffs[37] = 336;   // 0.020507 * 16384
    coeffs[38] = 360;   // 0.021956 * 16384
    coeffs[39] = 309;   // 0.018880 * 16384
    coeffs[40] = 215;   // 0.013124 * 16384
    coeffs[41] = 107;   // 0.006529 * 16384
    coeffs[42] = 10;    // 0.000602 * 16384
    coeffs[43] = -60;   // -0.003686 * 16384
    coeffs[44] = -98;   // -0.005959 * 16384
    coeffs[45] = -104;  // -0.006354 * 16384
    coeffs[46] = -88;   // -0.005364 * 16384
    coeffs[47] = -60;   // -0.003631 * 16384
    coeffs[48] = -29;   // -0.001766 * 16384
    coeffs[49] = -4;    // -0.000219 * 16384
    coeffs[50] = 13;    // 0.000778 * 16384
    coeffs[51] = 20;    // 0.001200 * 16384
    coeffs[52] = 19;    // 0.001169 * 16384
    coeffs[53] = 14;    // 0.000877 * 16384
    coeffs[54] = 8;     // 0.000511 * 16384
    coeffs[55] = 3;     // 0.000206 * 16384
    coeffs[56] = 0;     // 0.000024 * 16384

    end

    // Dãy mẫu đầu vào
    reg signed [15:0] x_reg [0:56];

    // Biến dùng trong xử lý
    integer i;
    reg signed [31:0] acc;

    always @(posedge clk) begin
        // Dịch dữ liệu
        for (i = 56; i > 0; i = i - 1)
            x_reg[i] <= x_reg[i - 1];
        x_reg[0] <= data_in;

        // Tính tích chập
        acc = 0;
        for (i = 0; i < 57; i = i + 1)
            acc = acc + x_reg[i] * coeffs[i];

        // Chia lại độ lớn (chuẩn Q1.14)
        data_out <= acc >>> 14;
    end

endmodule
